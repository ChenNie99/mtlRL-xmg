module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 ;
  assign n598 = x64 ^ x0 ^ 1'b0 ;
  assign n130 = x0 & x64 ;
  assign n129 = x65 ^ x1 ^ 1'b0 ;
  assign n131 = n130 ^ n129 ^ 1'b0 ;
  assign n133 = x1 & x65 ;
  assign n134 = n129 & n130 ;
  assign n135 = n133 | n134 ;
  assign n132 = x66 ^ x2 ^ 1'b0 ;
  assign n136 = n135 ^ n132 ^ 1'b0 ;
  assign n138 = x2 & x66 ;
  assign n139 = n132 & n135 ;
  assign n140 = n138 | n139 ;
  assign n137 = x67 ^ x3 ^ 1'b0 ;
  assign n141 = n140 ^ n137 ^ 1'b0 ;
  assign n143 = x3 & x67 ;
  assign n144 = n137 & n138 ;
  assign n145 = n143 | n144 ;
  assign n146 = n132 & n137 ;
  assign n147 = n135 & n146 ;
  assign n148 = n145 | n147 ;
  assign n142 = x68 ^ x4 ^ 1'b0 ;
  assign n149 = n148 ^ n142 ^ 1'b0 ;
  assign n151 = x4 & x68 ;
  assign n152 = n142 & n148 ;
  assign n153 = n151 | n152 ;
  assign n150 = x69 ^ x5 ^ 1'b0 ;
  assign n154 = n153 ^ n150 ^ 1'b0 ;
  assign n156 = x5 & x69 ;
  assign n157 = n150 & n151 ;
  assign n158 = n156 | n157 ;
  assign n159 = n142 & n150 ;
  assign n160 = n148 & n159 ;
  assign n161 = n158 | n160 ;
  assign n155 = x70 ^ x6 ^ 1'b0 ;
  assign n162 = n161 ^ n155 ^ 1'b0 ;
  assign n164 = x6 & x70 ;
  assign n165 = n155 & n161 ;
  assign n166 = n164 | n165 ;
  assign n163 = x71 ^ x7 ^ 1'b0 ;
  assign n167 = n166 ^ n163 ^ 1'b0 ;
  assign n169 = x7 & x71 ;
  assign n170 = n163 & n164 ;
  assign n171 = n169 | n170 ;
  assign n172 = n155 & n163 ;
  assign n173 = n158 & n172 ;
  assign n174 = n171 | n173 ;
  assign n175 = n159 & n172 ;
  assign n176 = n148 & n175 ;
  assign n177 = n174 | n176 ;
  assign n168 = x72 ^ x8 ^ 1'b0 ;
  assign n178 = n177 ^ n168 ^ 1'b0 ;
  assign n180 = x8 & x72 ;
  assign n181 = n168 & n177 ;
  assign n182 = n180 | n181 ;
  assign n179 = x73 ^ x9 ^ 1'b0 ;
  assign n183 = n182 ^ n179 ^ 1'b0 ;
  assign n185 = x9 & x73 ;
  assign n186 = n179 & n180 ;
  assign n187 = n185 | n186 ;
  assign n188 = n168 & n179 ;
  assign n189 = n177 & n188 ;
  assign n190 = n187 | n189 ;
  assign n184 = x74 ^ x10 ^ 1'b0 ;
  assign n191 = n190 ^ n184 ^ 1'b0 ;
  assign n193 = x10 & x74 ;
  assign n194 = n184 & n190 ;
  assign n195 = n193 | n194 ;
  assign n192 = x75 ^ x11 ^ 1'b0 ;
  assign n196 = n195 ^ n192 ^ 1'b0 ;
  assign n198 = x11 & x75 ;
  assign n199 = n192 & n193 ;
  assign n200 = n198 | n199 ;
  assign n201 = n184 & n192 ;
  assign n202 = n187 & n201 ;
  assign n203 = n200 | n202 ;
  assign n204 = n188 & n201 ;
  assign n205 = n177 & n204 ;
  assign n206 = n203 | n205 ;
  assign n197 = x76 ^ x12 ^ 1'b0 ;
  assign n207 = n206 ^ n197 ^ 1'b0 ;
  assign n209 = x12 & x76 ;
  assign n210 = n197 & n206 ;
  assign n211 = n209 | n210 ;
  assign n208 = x77 ^ x13 ^ 1'b0 ;
  assign n212 = n211 ^ n208 ^ 1'b0 ;
  assign n214 = x13 & x77 ;
  assign n215 = n208 & n209 ;
  assign n216 = n214 | n215 ;
  assign n217 = n197 & n208 ;
  assign n218 = n206 & n217 ;
  assign n219 = n216 | n218 ;
  assign n213 = x78 ^ x14 ^ 1'b0 ;
  assign n220 = n219 ^ n213 ^ 1'b0 ;
  assign n222 = x14 & x78 ;
  assign n223 = n213 & n219 ;
  assign n224 = n222 | n223 ;
  assign n221 = x79 ^ x15 ^ 1'b0 ;
  assign n225 = n224 ^ n221 ^ 1'b0 ;
  assign n227 = x15 & x79 ;
  assign n228 = n221 & n222 ;
  assign n229 = n227 | n228 ;
  assign n230 = n213 & n221 ;
  assign n231 = n216 & n230 ;
  assign n232 = n229 | n231 ;
  assign n233 = n217 & n230 ;
  assign n234 = n203 & n233 ;
  assign n235 = n232 | n234 ;
  assign n236 = n204 & n233 ;
  assign n237 = n177 & n236 ;
  assign n238 = n235 | n237 ;
  assign n226 = x80 ^ x16 ^ 1'b0 ;
  assign n239 = n238 ^ n226 ^ 1'b0 ;
  assign n241 = x16 & x80 ;
  assign n242 = n226 & n238 ;
  assign n243 = n241 | n242 ;
  assign n240 = x81 ^ x17 ^ 1'b0 ;
  assign n244 = n243 ^ n240 ^ 1'b0 ;
  assign n246 = x17 & x81 ;
  assign n247 = n240 & n241 ;
  assign n248 = n246 | n247 ;
  assign n249 = n226 & n240 ;
  assign n250 = n238 & n249 ;
  assign n251 = n248 | n250 ;
  assign n245 = x82 ^ x18 ^ 1'b0 ;
  assign n252 = n251 ^ n245 ^ 1'b0 ;
  assign n254 = x18 & x82 ;
  assign n255 = n245 & n251 ;
  assign n256 = n254 | n255 ;
  assign n253 = x83 ^ x19 ^ 1'b0 ;
  assign n257 = n256 ^ n253 ^ 1'b0 ;
  assign n259 = x19 & x83 ;
  assign n260 = n253 & n254 ;
  assign n261 = n259 | n260 ;
  assign n262 = n245 & n253 ;
  assign n263 = n248 & n262 ;
  assign n264 = n261 | n263 ;
  assign n265 = n249 & n262 ;
  assign n266 = n238 & n265 ;
  assign n267 = n264 | n266 ;
  assign n258 = x84 ^ x20 ^ 1'b0 ;
  assign n268 = n267 ^ n258 ^ 1'b0 ;
  assign n270 = x20 & x84 ;
  assign n271 = n258 & n267 ;
  assign n272 = n270 | n271 ;
  assign n269 = x85 ^ x21 ^ 1'b0 ;
  assign n273 = n272 ^ n269 ^ 1'b0 ;
  assign n275 = x21 & x85 ;
  assign n276 = n269 & n270 ;
  assign n277 = n275 | n276 ;
  assign n278 = n258 & n269 ;
  assign n279 = n267 & n278 ;
  assign n280 = n277 | n279 ;
  assign n274 = x86 ^ x22 ^ 1'b0 ;
  assign n281 = n280 ^ n274 ^ 1'b0 ;
  assign n283 = x22 & x86 ;
  assign n284 = n274 & n280 ;
  assign n285 = n283 | n284 ;
  assign n282 = x87 ^ x23 ^ 1'b0 ;
  assign n286 = n285 ^ n282 ^ 1'b0 ;
  assign n288 = x23 & x87 ;
  assign n289 = n282 & n283 ;
  assign n290 = n288 | n289 ;
  assign n291 = n274 & n282 ;
  assign n292 = n277 & n291 ;
  assign n293 = n290 | n292 ;
  assign n294 = n278 & n291 ;
  assign n295 = n264 & n294 ;
  assign n296 = n293 | n295 ;
  assign n297 = n265 & n294 ;
  assign n298 = n238 & n297 ;
  assign n299 = n296 | n298 ;
  assign n287 = x88 ^ x24 ^ 1'b0 ;
  assign n300 = n299 ^ n287 ^ 1'b0 ;
  assign n302 = x24 & x88 ;
  assign n303 = n287 & n299 ;
  assign n304 = n302 | n303 ;
  assign n301 = x89 ^ x25 ^ 1'b0 ;
  assign n305 = n304 ^ n301 ^ 1'b0 ;
  assign n307 = x25 & x89 ;
  assign n308 = n301 & n302 ;
  assign n309 = n307 | n308 ;
  assign n310 = n287 & n301 ;
  assign n311 = n299 & n310 ;
  assign n312 = n309 | n311 ;
  assign n306 = x90 ^ x26 ^ 1'b0 ;
  assign n313 = n312 ^ n306 ^ 1'b0 ;
  assign n315 = x26 & x90 ;
  assign n316 = n306 & n312 ;
  assign n317 = n315 | n316 ;
  assign n314 = x91 ^ x27 ^ 1'b0 ;
  assign n318 = n317 ^ n314 ^ 1'b0 ;
  assign n320 = x27 & x91 ;
  assign n321 = n314 & n315 ;
  assign n322 = n320 | n321 ;
  assign n323 = n306 & n314 ;
  assign n324 = n309 & n323 ;
  assign n325 = n322 | n324 ;
  assign n326 = n310 & n323 ;
  assign n327 = n299 & n326 ;
  assign n328 = n325 | n327 ;
  assign n319 = x92 ^ x28 ^ 1'b0 ;
  assign n329 = n328 ^ n319 ^ 1'b0 ;
  assign n331 = x28 & x92 ;
  assign n332 = n319 & n328 ;
  assign n333 = n331 | n332 ;
  assign n330 = x93 ^ x29 ^ 1'b0 ;
  assign n334 = n333 ^ n330 ^ 1'b0 ;
  assign n336 = x29 & x93 ;
  assign n337 = n330 & n331 ;
  assign n338 = n336 | n337 ;
  assign n339 = n319 & n330 ;
  assign n340 = n328 & n339 ;
  assign n341 = n338 | n340 ;
  assign n335 = x94 ^ x30 ^ 1'b0 ;
  assign n342 = n341 ^ n335 ^ 1'b0 ;
  assign n344 = x30 & x94 ;
  assign n345 = n335 & n341 ;
  assign n346 = n344 | n345 ;
  assign n343 = x95 ^ x31 ^ 1'b0 ;
  assign n347 = n346 ^ n343 ^ 1'b0 ;
  assign n349 = x31 & x95 ;
  assign n350 = n343 & n344 ;
  assign n351 = n349 | n350 ;
  assign n352 = n335 & n343 ;
  assign n353 = n338 & n352 ;
  assign n354 = n351 | n353 ;
  assign n355 = n339 & n352 ;
  assign n356 = n325 & n355 ;
  assign n357 = n354 | n356 ;
  assign n358 = n326 & n355 ;
  assign n359 = n296 & n358 ;
  assign n360 = n357 | n359 ;
  assign n361 = n297 & n358 ;
  assign n362 = n238 & n361 ;
  assign n363 = n360 | n362 ;
  assign n348 = x96 ^ x32 ^ 1'b0 ;
  assign n364 = n363 ^ n348 ^ 1'b0 ;
  assign n366 = x32 & x96 ;
  assign n367 = n348 & n363 ;
  assign n368 = n366 | n367 ;
  assign n365 = x97 ^ x33 ^ 1'b0 ;
  assign n369 = n368 ^ n365 ^ 1'b0 ;
  assign n371 = x33 & x97 ;
  assign n372 = n365 & n366 ;
  assign n373 = n371 | n372 ;
  assign n374 = n348 & n365 ;
  assign n375 = n363 & n374 ;
  assign n376 = n373 | n375 ;
  assign n370 = x98 ^ x34 ^ 1'b0 ;
  assign n377 = n376 ^ n370 ^ 1'b0 ;
  assign n379 = x34 & x98 ;
  assign n380 = n370 & n376 ;
  assign n381 = n379 | n380 ;
  assign n378 = x99 ^ x35 ^ 1'b0 ;
  assign n382 = n381 ^ n378 ^ 1'b0 ;
  assign n384 = x35 & x99 ;
  assign n385 = n378 & n379 ;
  assign n386 = n384 | n385 ;
  assign n387 = n370 & n378 ;
  assign n388 = n373 & n387 ;
  assign n389 = n386 | n388 ;
  assign n390 = n374 & n387 ;
  assign n391 = n363 & n390 ;
  assign n392 = n389 | n391 ;
  assign n383 = x100 ^ x36 ^ 1'b0 ;
  assign n393 = n392 ^ n383 ^ 1'b0 ;
  assign n395 = x36 & x100 ;
  assign n396 = n383 & n392 ;
  assign n397 = n395 | n396 ;
  assign n394 = x101 ^ x37 ^ 1'b0 ;
  assign n398 = n397 ^ n394 ^ 1'b0 ;
  assign n400 = n394 & n395 ;
  assign n401 = x37 & x101 ;
  assign n402 = n400 | n401 ;
  assign n403 = n383 & n394 ;
  assign n404 = n392 & n403 ;
  assign n405 = n402 | n404 ;
  assign n399 = x102 ^ x38 ^ 1'b0 ;
  assign n406 = n405 ^ n399 ^ 1'b0 ;
  assign n408 = x38 & x102 ;
  assign n409 = n399 & n405 ;
  assign n410 = n408 | n409 ;
  assign n407 = x103 ^ x39 ^ 1'b0 ;
  assign n411 = n410 ^ n407 ^ 1'b0 ;
  assign n413 = x39 & x103 ;
  assign n414 = n407 & n408 ;
  assign n415 = n413 | n414 ;
  assign n416 = n399 & n407 ;
  assign n417 = n402 & n416 ;
  assign n418 = n415 | n417 ;
  assign n419 = n403 & n416 ;
  assign n420 = n389 & n419 ;
  assign n421 = n418 | n420 ;
  assign n422 = n390 & n419 ;
  assign n423 = n363 & n422 ;
  assign n424 = n421 | n423 ;
  assign n412 = x104 ^ x40 ^ 1'b0 ;
  assign n425 = n424 ^ n412 ^ 1'b0 ;
  assign n427 = x40 & x104 ;
  assign n428 = n412 & n424 ;
  assign n429 = n427 | n428 ;
  assign n426 = x105 ^ x41 ^ 1'b0 ;
  assign n430 = n429 ^ n426 ^ 1'b0 ;
  assign n432 = n426 & n427 ;
  assign n433 = x41 & x105 ;
  assign n434 = n432 | n433 ;
  assign n435 = n412 & n426 ;
  assign n436 = n424 & n435 ;
  assign n437 = n434 | n436 ;
  assign n431 = x106 ^ x42 ^ 1'b0 ;
  assign n438 = n437 ^ n431 ^ 1'b0 ;
  assign n440 = x42 & x106 ;
  assign n441 = n431 & n437 ;
  assign n442 = n440 | n441 ;
  assign n439 = x107 ^ x43 ^ 1'b0 ;
  assign n443 = n442 ^ n439 ^ 1'b0 ;
  assign n445 = x43 & x107 ;
  assign n446 = n439 & n440 ;
  assign n447 = n445 | n446 ;
  assign n448 = n431 & n439 ;
  assign n449 = n434 & n448 ;
  assign n450 = n447 | n449 ;
  assign n451 = n435 & n448 ;
  assign n452 = n424 & n451 ;
  assign n453 = n450 | n452 ;
  assign n444 = x108 ^ x44 ^ 1'b0 ;
  assign n454 = n453 ^ n444 ^ 1'b0 ;
  assign n456 = x44 & x108 ;
  assign n457 = n444 & n453 ;
  assign n458 = n456 | n457 ;
  assign n455 = x109 ^ x45 ^ 1'b0 ;
  assign n459 = n458 ^ n455 ^ 1'b0 ;
  assign n461 = x45 & x109 ;
  assign n462 = n455 & n456 ;
  assign n463 = n461 | n462 ;
  assign n464 = n444 & n455 ;
  assign n465 = n453 & n464 ;
  assign n466 = n463 | n465 ;
  assign n460 = x110 ^ x46 ^ 1'b0 ;
  assign n467 = n466 ^ n460 ^ 1'b0 ;
  assign n469 = x46 & x110 ;
  assign n470 = n460 & n466 ;
  assign n471 = n469 | n470 ;
  assign n468 = x111 ^ x47 ^ 1'b0 ;
  assign n472 = n471 ^ n468 ^ 1'b0 ;
  assign n474 = x47 & x111 ;
  assign n475 = n468 & n469 ;
  assign n476 = n474 | n475 ;
  assign n477 = n460 & n468 ;
  assign n478 = n463 & n477 ;
  assign n479 = n476 | n478 ;
  assign n480 = n464 & n477 ;
  assign n481 = n450 & n480 ;
  assign n482 = n479 | n481 ;
  assign n483 = n451 & n480 ;
  assign n484 = n421 & n483 ;
  assign n485 = n482 | n484 ;
  assign n486 = n422 & n483 ;
  assign n487 = n363 & n486 ;
  assign n488 = n485 | n487 ;
  assign n473 = x112 ^ x48 ^ 1'b0 ;
  assign n489 = n488 ^ n473 ^ 1'b0 ;
  assign n491 = x48 & x112 ;
  assign n492 = n473 & n488 ;
  assign n493 = n491 | n492 ;
  assign n490 = x113 ^ x49 ^ 1'b0 ;
  assign n494 = n493 ^ n490 ^ 1'b0 ;
  assign n496 = x49 & x113 ;
  assign n497 = n490 & n491 ;
  assign n498 = n496 | n497 ;
  assign n499 = n473 & n490 ;
  assign n500 = n488 & n499 ;
  assign n501 = n498 | n500 ;
  assign n495 = x114 ^ x50 ^ 1'b0 ;
  assign n502 = n501 ^ n495 ^ 1'b0 ;
  assign n504 = x50 & x114 ;
  assign n505 = n495 & n501 ;
  assign n506 = n504 | n505 ;
  assign n503 = x115 ^ x51 ^ 1'b0 ;
  assign n507 = n506 ^ n503 ^ 1'b0 ;
  assign n509 = x51 & x115 ;
  assign n510 = n503 & n504 ;
  assign n511 = n509 | n510 ;
  assign n512 = n495 & n503 ;
  assign n513 = n498 & n512 ;
  assign n514 = n511 | n513 ;
  assign n515 = n499 & n512 ;
  assign n516 = n488 & n515 ;
  assign n517 = n514 | n516 ;
  assign n508 = x116 ^ x52 ^ 1'b0 ;
  assign n518 = n517 ^ n508 ^ 1'b0 ;
  assign n520 = x52 & x116 ;
  assign n521 = n508 & n517 ;
  assign n522 = n520 | n521 ;
  assign n519 = x117 ^ x53 ^ 1'b0 ;
  assign n523 = n522 ^ n519 ^ 1'b0 ;
  assign n525 = x53 & x117 ;
  assign n526 = n519 & n520 ;
  assign n527 = n525 | n526 ;
  assign n528 = n508 & n519 ;
  assign n529 = n517 & n528 ;
  assign n530 = n527 | n529 ;
  assign n524 = x118 ^ x54 ^ 1'b0 ;
  assign n531 = n530 ^ n524 ^ 1'b0 ;
  assign n533 = x54 & x118 ;
  assign n534 = n524 & n530 ;
  assign n535 = n533 | n534 ;
  assign n532 = x119 ^ x55 ^ 1'b0 ;
  assign n536 = n535 ^ n532 ^ 1'b0 ;
  assign n538 = x55 & x119 ;
  assign n539 = n532 & n533 ;
  assign n540 = n538 | n539 ;
  assign n541 = n524 & n532 ;
  assign n542 = n527 & n541 ;
  assign n543 = n540 | n542 ;
  assign n544 = n528 & n541 ;
  assign n545 = n514 & n544 ;
  assign n546 = n543 | n545 ;
  assign n547 = n515 & n544 ;
  assign n548 = n488 & n547 ;
  assign n549 = n546 | n548 ;
  assign n537 = x120 ^ x56 ^ 1'b0 ;
  assign n550 = n549 ^ n537 ^ 1'b0 ;
  assign n552 = x56 & x120 ;
  assign n553 = n537 & n549 ;
  assign n554 = n552 | n553 ;
  assign n551 = x121 ^ x57 ^ 1'b0 ;
  assign n555 = n554 ^ n551 ^ 1'b0 ;
  assign n557 = n551 & n552 ;
  assign n558 = x57 & x121 ;
  assign n559 = n557 | n558 ;
  assign n560 = n537 & n551 ;
  assign n561 = n549 & n560 ;
  assign n562 = n559 | n561 ;
  assign n556 = x122 ^ x58 ^ 1'b0 ;
  assign n563 = n562 ^ n556 ^ 1'b0 ;
  assign n565 = x58 & x122 ;
  assign n566 = n556 & n562 ;
  assign n567 = n565 | n566 ;
  assign n564 = x123 ^ x59 ^ 1'b0 ;
  assign n568 = n567 ^ n564 ^ 1'b0 ;
  assign n570 = n564 & n565 ;
  assign n571 = x59 & x123 ;
  assign n572 = n570 | n571 ;
  assign n573 = n556 & n564 ;
  assign n574 = n559 & n573 ;
  assign n575 = n572 | n574 ;
  assign n576 = n560 & n573 ;
  assign n577 = n549 & n576 ;
  assign n578 = n575 | n577 ;
  assign n569 = x124 ^ x60 ^ 1'b0 ;
  assign n579 = n578 ^ n569 ^ 1'b0 ;
  assign n581 = x60 & x124 ;
  assign n582 = n569 & n578 ;
  assign n583 = n581 | n582 ;
  assign n580 = x125 ^ x61 ^ 1'b0 ;
  assign n584 = n583 ^ n580 ^ 1'b0 ;
  assign n586 = n580 & n581 ;
  assign n587 = x61 & x125 ;
  assign n588 = n586 | n587 ;
  assign n589 = n569 & n580 ;
  assign n590 = n578 & n589 ;
  assign n591 = n588 | n590 ;
  assign n585 = x126 ^ x62 ^ 1'b0 ;
  assign n592 = n591 ^ n585 ^ 1'b0 ;
  assign n594 = x62 & x126 ;
  assign n595 = n585 & n591 ;
  assign n596 = n594 | n595 ;
  assign n593 = x127 ^ x63 ^ 1'b0 ;
  assign n597 = n596 ^ n593 ^ 1'b0 ;
  assign y0 = n598 ;
  assign y1 = n131 ;
  assign y2 = n136 ;
  assign y3 = n141 ;
  assign y4 = n149 ;
  assign y5 = n154 ;
  assign y6 = n162 ;
  assign y7 = n167 ;
  assign y8 = n178 ;
  assign y9 = n183 ;
  assign y10 = n191 ;
  assign y11 = n196 ;
  assign y12 = n207 ;
  assign y13 = n212 ;
  assign y14 = n220 ;
  assign y15 = n225 ;
  assign y16 = n239 ;
  assign y17 = n244 ;
  assign y18 = n252 ;
  assign y19 = n257 ;
  assign y20 = n268 ;
  assign y21 = n273 ;
  assign y22 = n281 ;
  assign y23 = n286 ;
  assign y24 = n300 ;
  assign y25 = n305 ;
  assign y26 = n313 ;
  assign y27 = n318 ;
  assign y28 = n329 ;
  assign y29 = n334 ;
  assign y30 = n342 ;
  assign y31 = n347 ;
  assign y32 = n364 ;
  assign y33 = n369 ;
  assign y34 = n377 ;
  assign y35 = n382 ;
  assign y36 = n393 ;
  assign y37 = n398 ;
  assign y38 = n406 ;
  assign y39 = n411 ;
  assign y40 = n425 ;
  assign y41 = n430 ;
  assign y42 = n438 ;
  assign y43 = n443 ;
  assign y44 = n454 ;
  assign y45 = n459 ;
  assign y46 = n467 ;
  assign y47 = n472 ;
  assign y48 = n489 ;
  assign y49 = n494 ;
  assign y50 = n502 ;
  assign y51 = n507 ;
  assign y52 = n518 ;
  assign y53 = n523 ;
  assign y54 = n531 ;
  assign y55 = n536 ;
  assign y56 = n550 ;
  assign y57 = n555 ;
  assign y58 = n563 ;
  assign y59 = n568 ;
  assign y60 = n579 ;
  assign y61 = n584 ;
  assign y62 = n592 ;
  assign y63 = n597 ;
endmodule
