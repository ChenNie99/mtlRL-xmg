module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 ;
  assign n47 = x16 ^ x15 ^ x13 ;
  assign n48 = n47 ^ x14 ^ 1'b0 ;
  assign n45 = x12 ^ x10 ^ x8 ;
  assign n46 = n45 ^ x9 ^ 1'b0 ;
  assign n49 = n48 ^ n46 ^ 1'b0 ;
  assign n43 = x40 ^ x36 ^ x0 ;
  assign n44 = n43 ^ x4 ^ 1'b0 ;
  assign n50 = n49 ^ n44 ^ 1'b0 ;
  assign n42 = x26 & x35 ;
  assign n51 = n50 ^ n42 ^ 1'b0 ;
  assign n58 = x32 & x35 ;
  assign n56 = x24 ^ x19 ^ x10 ;
  assign n57 = n56 ^ x15 ^ 1'b0 ;
  assign n59 = n58 ^ n57 ^ 1'b0 ;
  assign n54 = x33 ^ x22 ^ x0 ;
  assign n55 = n54 ^ x11 ^ 1'b0 ;
  assign n60 = n59 ^ n55 ^ 1'b0 ;
  assign n52 = x40 ^ x3 ^ x1 ;
  assign n53 = n52 ^ x2 ^ 1'b0 ;
  assign n61 = n60 ^ n53 ^ 1'b0 ;
  assign n65 = x25 ^ x24 ^ x21 ;
  assign n66 = n65 ^ x23 ^ 1'b0 ;
  assign n64 = x29 & x35 ;
  assign n67 = n66 ^ n64 ^ 1'b0 ;
  assign n68 = n67 ^ n48 ^ 1'b0 ;
  assign n62 = x39 ^ x33 ^ x3 ;
  assign n63 = n62 ^ x7 ^ 1'b0 ;
  assign n69 = n68 ^ n63 ^ 1'b0 ;
  assign n74 = x28 & x35 ;
  assign n72 = x38 ^ x22 ^ x2 ;
  assign n73 = n72 ^ x6 ^ 1'b0 ;
  assign n75 = n74 ^ n73 ^ 1'b0 ;
  assign n76 = n75 ^ n46 ^ 1'b0 ;
  assign n70 = x20 ^ x19 ^ x17 ;
  assign n71 = n70 ^ x18 ^ 1'b0 ;
  assign n77 = n76 ^ n71 ^ 1'b0 ;
  assign n78 = ( n51 & n69 ) | ( n51 & n77 ) | ( n69 & n77 ) ;
  assign n85 = n69 ^ n51 ^ 1'b0 ;
  assign n86 = ( n77 & ~n78 ) | ( n77 & n85 ) | ( ~n78 & n85 ) ;
  assign n81 = x27 & x35 ;
  assign n82 = n81 ^ n71 ^ 1'b0 ;
  assign n83 = n82 ^ n66 ^ 1'b0 ;
  assign n79 = x37 ^ x11 ^ x1 ;
  assign n80 = n79 ^ x5 ^ 1'b0 ;
  assign n84 = n83 ^ n80 ^ 1'b0 ;
  assign n87 = n86 ^ n84 ^ 1'b0 ;
  assign n88 = ~n78 & n87 ;
  assign n89 = n61 & n88 ;
  assign n93 = x39 ^ x38 ^ x36 ;
  assign n94 = n93 ^ x37 ^ 1'b0 ;
  assign n95 = n94 ^ n55 ^ 1'b0 ;
  assign n91 = x21 ^ x17 ^ x8 ;
  assign n92 = n91 ^ x13 ^ 1'b0 ;
  assign n96 = n95 ^ n92 ^ 1'b0 ;
  assign n90 = x30 & x35 ;
  assign n97 = n96 ^ n90 ^ 1'b0 ;
  assign n101 = x7 ^ x6 ^ x4 ;
  assign n102 = n101 ^ x5 ^ 1'b0 ;
  assign n103 = n102 ^ n53 ^ 1'b0 ;
  assign n99 = x23 ^ x18 ^ x9 ;
  assign n100 = n99 ^ x14 ^ 1'b0 ;
  assign n104 = n103 ^ n100 ^ 1'b0 ;
  assign n98 = x31 & x35 ;
  assign n105 = n104 ^ n98 ^ 1'b0 ;
  assign n106 = n97 & ~n105 ;
  assign n109 = x34 & x35 ;
  assign n107 = x25 ^ x20 ^ x12 ;
  assign n108 = n107 ^ x16 ^ 1'b0 ;
  assign n110 = n109 ^ n108 ^ 1'b0 ;
  assign n111 = n110 ^ n94 ^ 1'b0 ;
  assign n112 = n111 ^ n102 ^ 1'b0 ;
  assign n113 = ( n61 & ~n106 ) | ( n61 & n112 ) | ( ~n106 & n112 ) ;
  assign n114 = n89 & ~n113 ;
  assign n115 = n51 & n114 ;
  assign n116 = n115 ^ x0 ^ 1'b0 ;
  assign n117 = n84 & n114 ;
  assign n118 = n117 ^ x11 ^ 1'b0 ;
  assign n119 = n77 & n114 ;
  assign n120 = n119 ^ x22 ^ 1'b0 ;
  assign n121 = n69 & n114 ;
  assign n122 = n121 ^ x33 ^ 1'b0 ;
  assign n123 = ~n61 & n88 ;
  assign n124 = ( n61 & n106 ) | ( n61 & n112 ) | ( n106 & n112 ) ;
  assign n125 = n123 & n124 ;
  assign n126 = n51 & n125 ;
  assign n127 = n126 ^ x36 ^ 1'b0 ;
  assign n128 = n84 & n125 ;
  assign n129 = n128 ^ x37 ^ 1'b0 ;
  assign n130 = n77 & n125 ;
  assign n131 = n130 ^ x38 ^ 1'b0 ;
  assign n132 = n69 & n125 ;
  assign n133 = n132 ^ x39 ^ 1'b0 ;
  assign n134 = ~n97 & n105 ;
  assign n135 = ~n112 & n134 ;
  assign n136 = ( n61 & n88 ) | ( n61 & n112 ) | ( n88 & n112 ) ;
  assign n137 = n135 & n136 ;
  assign n138 = n51 & n137 ;
  assign n139 = n138 ^ x40 ^ 1'b0 ;
  assign n140 = n84 & n137 ;
  assign n141 = n140 ^ x1 ^ 1'b0 ;
  assign n142 = n77 & n137 ;
  assign n143 = n142 ^ x2 ^ 1'b0 ;
  assign n144 = n69 & n137 ;
  assign n145 = n144 ^ x3 ^ 1'b0 ;
  assign n146 = n112 & n134 ;
  assign n147 = ( n61 & ~n88 ) | ( n61 & n112 ) | ( ~n88 & n112 ) ;
  assign n148 = n146 & ~n147 ;
  assign n149 = n51 & n148 ;
  assign n150 = n149 ^ x4 ^ 1'b0 ;
  assign n151 = n84 & n148 ;
  assign n152 = n151 ^ x5 ^ 1'b0 ;
  assign n153 = n77 & n148 ;
  assign n154 = n153 ^ x6 ^ 1'b0 ;
  assign n155 = n69 & n148 ;
  assign n156 = n155 ^ x7 ^ 1'b0 ;
  assign n157 = ( n97 & n105 ) | ( n97 & n112 ) | ( n105 & n112 ) ;
  assign n158 = n105 ^ n97 ^ 1'b0 ;
  assign n159 = ( n112 & ~n157 ) | ( n112 & n158 ) | ( ~n157 & n158 ) ;
  assign n160 = n159 ^ n61 ^ 1'b0 ;
  assign n161 = ~n157 & n160 ;
  assign n162 = n77 & n161 ;
  assign n163 = n51 & ~n84 ;
  assign n164 = ( n69 & n77 ) | ( n69 & ~n163 ) | ( n77 & ~n163 ) ;
  assign n165 = n162 & ~n164 ;
  assign n166 = n97 & n165 ;
  assign n167 = n166 ^ x8 ^ 1'b0 ;
  assign n168 = n105 & n165 ;
  assign n169 = n168 ^ x9 ^ 1'b0 ;
  assign n170 = n61 & n165 ;
  assign n171 = n170 ^ x10 ^ 1'b0 ;
  assign n172 = n112 & n165 ;
  assign n173 = n172 ^ x12 ^ 1'b0 ;
  assign n174 = ~n77 & n161 ;
  assign n175 = ( n69 & n77 ) | ( n69 & n163 ) | ( n77 & n163 ) ;
  assign n176 = n174 & n175 ;
  assign n177 = n97 & n176 ;
  assign n178 = n177 ^ x13 ^ 1'b0 ;
  assign n179 = n105 & n176 ;
  assign n180 = n179 ^ x14 ^ 1'b0 ;
  assign n181 = n61 & n176 ;
  assign n182 = n181 ^ x15 ^ 1'b0 ;
  assign n183 = n112 & n176 ;
  assign n184 = n183 ^ x16 ^ 1'b0 ;
  assign n185 = ~n51 & n84 ;
  assign n186 = ( n69 & n77 ) | ( n69 & ~n185 ) | ( n77 & ~n185 ) ;
  assign n187 = n162 & ~n186 ;
  assign n188 = n97 & n187 ;
  assign n189 = n188 ^ x17 ^ 1'b0 ;
  assign n190 = n105 & n187 ;
  assign n191 = n190 ^ x18 ^ 1'b0 ;
  assign n192 = n61 & n187 ;
  assign n193 = n192 ^ x19 ^ 1'b0 ;
  assign n194 = n112 & n187 ;
  assign n195 = n194 ^ x20 ^ 1'b0 ;
  assign n196 = ( n69 & n77 ) | ( n69 & n185 ) | ( n77 & n185 ) ;
  assign n197 = n174 & n196 ;
  assign n198 = n97 & n197 ;
  assign n199 = n198 ^ x21 ^ 1'b0 ;
  assign n200 = n105 & n197 ;
  assign n201 = n200 ^ x23 ^ 1'b0 ;
  assign n202 = n61 & n197 ;
  assign n203 = n202 ^ x24 ^ 1'b0 ;
  assign n204 = n112 & n197 ;
  assign n205 = n204 ^ x25 ^ 1'b0 ;
  assign y0 = ~n116 ;
  assign y1 = ~n118 ;
  assign y2 = ~n120 ;
  assign y3 = ~n122 ;
  assign y4 = ~n127 ;
  assign y5 = ~n129 ;
  assign y6 = ~n131 ;
  assign y7 = ~n133 ;
  assign y8 = ~n139 ;
  assign y9 = ~n141 ;
  assign y10 = ~n143 ;
  assign y11 = ~n145 ;
  assign y12 = ~n150 ;
  assign y13 = ~n152 ;
  assign y14 = ~n154 ;
  assign y15 = ~n156 ;
  assign y16 = ~n167 ;
  assign y17 = ~n169 ;
  assign y18 = ~n171 ;
  assign y19 = ~n173 ;
  assign y20 = ~n178 ;
  assign y21 = ~n180 ;
  assign y22 = ~n182 ;
  assign y23 = ~n184 ;
  assign y24 = ~n189 ;
  assign y25 = ~n191 ;
  assign y26 = ~n193 ;
  assign y27 = ~n195 ;
  assign y28 = ~n199 ;
  assign y29 = ~n201 ;
  assign y30 = ~n203 ;
  assign y31 = ~n205 ;
endmodule
