module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 ;
  assign n129 = x64 ^ x0 ^ 1'b0 ;
  assign n130 = x0 & x64 ;
  assign n131 = n130 ^ x65 ^ x1 ;
  assign n133 = x66 ^ x2 ^ 1'b0 ;
  assign n132 = ( x1 & x65 ) | ( x1 & n130 ) | ( x65 & n130 ) ;
  assign n134 = n133 ^ n132 ^ 1'b0 ;
  assign n136 = ( x2 & x66 ) | ( x2 & n132 ) | ( x66 & n132 ) ;
  assign n135 = x67 ^ x3 ^ 1'b0 ;
  assign n137 = n136 ^ n135 ^ 1'b0 ;
  assign n143 = x68 ^ x4 ^ 1'b0 ;
  assign n138 = x2 & x66 ;
  assign n139 = ( x3 & x67 ) | ( x3 & n138 ) | ( x67 & n138 ) ;
  assign n140 = n132 & ~n133 ;
  assign n141 = ( n132 & n135 ) | ( n132 & n140 ) | ( n135 & n140 ) ;
  assign n142 = ( n139 & ~n140 ) | ( n139 & n141 ) | ( ~n140 & n141 ) ;
  assign n144 = n143 ^ n142 ^ 1'b0 ;
  assign n146 = ( x4 & x68 ) | ( x4 & n142 ) | ( x68 & n142 ) ;
  assign n145 = x69 ^ x5 ^ 1'b0 ;
  assign n147 = n146 ^ n145 ^ 1'b0 ;
  assign n153 = x70 ^ x6 ^ 1'b0 ;
  assign n148 = x4 & x68 ;
  assign n149 = ( x5 & x69 ) | ( x5 & n148 ) | ( x69 & n148 ) ;
  assign n150 = n143 & n145 ;
  assign n151 = ( n142 & n149 ) | ( n142 & n150 ) | ( n149 & n150 ) ;
  assign n152 = n149 | n151 ;
  assign n154 = n153 ^ n152 ^ 1'b0 ;
  assign n156 = ( x6 & x70 ) | ( x6 & n152 ) | ( x70 & n152 ) ;
  assign n155 = x71 ^ x7 ^ 1'b0 ;
  assign n157 = n156 ^ n155 ^ 1'b0 ;
  assign n166 = x72 ^ x8 ^ 1'b0 ;
  assign n158 = x6 & x70 ;
  assign n159 = ( x7 & x71 ) | ( x7 & n158 ) | ( x71 & n158 ) ;
  assign n160 = n153 & n155 ;
  assign n161 = ( n149 & n159 ) | ( n149 & n160 ) | ( n159 & n160 ) ;
  assign n162 = n159 | n161 ;
  assign n163 = ~n142 & n150 ;
  assign n164 = ( n150 & n160 ) | ( n150 & n163 ) | ( n160 & n163 ) ;
  assign n165 = ( n162 & ~n163 ) | ( n162 & n164 ) | ( ~n163 & n164 ) ;
  assign n167 = n166 ^ n165 ^ 1'b0 ;
  assign n169 = ( x8 & x72 ) | ( x8 & n165 ) | ( x72 & n165 ) ;
  assign n168 = x73 ^ x9 ^ 1'b0 ;
  assign n170 = n169 ^ n168 ^ 1'b0 ;
  assign n176 = x74 ^ x10 ^ 1'b0 ;
  assign n171 = x8 & x72 ;
  assign n172 = ( x9 & x73 ) | ( x9 & n171 ) | ( x73 & n171 ) ;
  assign n173 = n166 & n168 ;
  assign n174 = ( n165 & n172 ) | ( n165 & n173 ) | ( n172 & n173 ) ;
  assign n175 = n172 | n174 ;
  assign n177 = n176 ^ n175 ^ 1'b0 ;
  assign n179 = ( x10 & x74 ) | ( x10 & n175 ) | ( x74 & n175 ) ;
  assign n178 = x75 ^ x11 ^ 1'b0 ;
  assign n180 = n179 ^ n178 ^ 1'b0 ;
  assign n190 = x76 ^ x12 ^ 1'b0 ;
  assign n181 = x10 & x74 ;
  assign n182 = ( x11 & x75 ) | ( x11 & n181 ) | ( x75 & n181 ) ;
  assign n183 = n176 & n178 ;
  assign n184 = ( n172 & n182 ) | ( n172 & n183 ) | ( n182 & n183 ) ;
  assign n185 = n182 | n184 ;
  assign n186 = ( n173 & n176 ) | ( n173 & ~n178 ) | ( n176 & ~n178 ) ;
  assign n187 = n178 & n186 ;
  assign n188 = ( n165 & n185 ) | ( n165 & n187 ) | ( n185 & n187 ) ;
  assign n189 = n185 | n188 ;
  assign n191 = n190 ^ n189 ^ 1'b0 ;
  assign n193 = ( x12 & x76 ) | ( x12 & n189 ) | ( x76 & n189 ) ;
  assign n192 = x77 ^ x13 ^ 1'b0 ;
  assign n194 = n193 ^ n192 ^ 1'b0 ;
  assign n200 = x78 ^ x14 ^ 1'b0 ;
  assign n195 = x12 & x76 ;
  assign n196 = ( x13 & x77 ) | ( x13 & n195 ) | ( x77 & n195 ) ;
  assign n197 = n190 & n192 ;
  assign n198 = ( n189 & n196 ) | ( n189 & n197 ) | ( n196 & n197 ) ;
  assign n199 = n196 | n198 ;
  assign n201 = n200 ^ n199 ^ 1'b0 ;
  assign n203 = ( x14 & x78 ) | ( x14 & n199 ) | ( x78 & n199 ) ;
  assign n202 = x79 ^ x15 ^ 1'b0 ;
  assign n204 = n203 ^ n202 ^ 1'b0 ;
  assign n217 = x80 ^ x16 ^ 1'b0 ;
  assign n205 = x14 & x78 ;
  assign n206 = ( x15 & x79 ) | ( x15 & n205 ) | ( x79 & n205 ) ;
  assign n207 = ( n196 & n200 ) | ( n196 & ~n202 ) | ( n200 & ~n202 ) ;
  assign n208 = n202 & n207 ;
  assign n209 = n206 | n208 ;
  assign n210 = ( n197 & n200 ) | ( n197 & ~n202 ) | ( n200 & ~n202 ) ;
  assign n211 = n202 & n210 ;
  assign n212 = ( n185 & n208 ) | ( n185 & n211 ) | ( n208 & n211 ) ;
  assign n213 = n209 | n212 ;
  assign n214 = ~n165 & n187 ;
  assign n215 = ( n187 & n211 ) | ( n187 & n214 ) | ( n211 & n214 ) ;
  assign n216 = ( n213 & ~n214 ) | ( n213 & n215 ) | ( ~n214 & n215 ) ;
  assign n218 = n217 ^ n216 ^ 1'b0 ;
  assign n220 = ( x16 & x80 ) | ( x16 & n216 ) | ( x80 & n216 ) ;
  assign n219 = x81 ^ x17 ^ 1'b0 ;
  assign n221 = n220 ^ n219 ^ 1'b0 ;
  assign n227 = x82 ^ x18 ^ 1'b0 ;
  assign n222 = x16 & x80 ;
  assign n223 = ( x17 & x81 ) | ( x17 & n222 ) | ( x81 & n222 ) ;
  assign n224 = n217 & n219 ;
  assign n225 = ( n216 & n223 ) | ( n216 & n224 ) | ( n223 & n224 ) ;
  assign n226 = n223 | n225 ;
  assign n228 = n227 ^ n226 ^ 1'b0 ;
  assign n230 = ( x18 & x82 ) | ( x18 & n226 ) | ( x82 & n226 ) ;
  assign n229 = x83 ^ x19 ^ 1'b0 ;
  assign n231 = n230 ^ n229 ^ 1'b0 ;
  assign n241 = x84 ^ x20 ^ 1'b0 ;
  assign n232 = x18 & x82 ;
  assign n233 = ( x19 & x83 ) | ( x19 & n232 ) | ( x83 & n232 ) ;
  assign n234 = n227 & n229 ;
  assign n235 = ( n223 & n233 ) | ( n223 & n234 ) | ( n233 & n234 ) ;
  assign n236 = n233 | n235 ;
  assign n237 = ( n224 & n227 ) | ( n224 & ~n229 ) | ( n227 & ~n229 ) ;
  assign n238 = n229 & n237 ;
  assign n239 = ( n216 & n236 ) | ( n216 & n238 ) | ( n236 & n238 ) ;
  assign n240 = n236 | n239 ;
  assign n242 = n241 ^ n240 ^ 1'b0 ;
  assign n244 = ( x20 & x84 ) | ( x20 & n240 ) | ( x84 & n240 ) ;
  assign n243 = x85 ^ x21 ^ 1'b0 ;
  assign n245 = n244 ^ n243 ^ 1'b0 ;
  assign n251 = x86 ^ x22 ^ 1'b0 ;
  assign n246 = x20 & x84 ;
  assign n247 = ( x21 & x85 ) | ( x21 & n246 ) | ( x85 & n246 ) ;
  assign n248 = n241 & n243 ;
  assign n249 = ( n240 & n247 ) | ( n240 & n248 ) | ( n247 & n248 ) ;
  assign n250 = n247 | n249 ;
  assign n252 = n251 ^ n250 ^ 1'b0 ;
  assign n254 = ( x22 & x86 ) | ( x22 & n250 ) | ( x86 & n250 ) ;
  assign n253 = x87 ^ x23 ^ 1'b0 ;
  assign n255 = n254 ^ n253 ^ 1'b0 ;
  assign n268 = x88 ^ x24 ^ 1'b0 ;
  assign n256 = x22 & x86 ;
  assign n257 = ( x23 & x87 ) | ( x23 & n256 ) | ( x87 & n256 ) ;
  assign n258 = ( n247 & n251 ) | ( n247 & ~n253 ) | ( n251 & ~n253 ) ;
  assign n259 = n253 & n258 ;
  assign n260 = n257 | n259 ;
  assign n261 = ( n248 & n251 ) | ( n248 & ~n253 ) | ( n251 & ~n253 ) ;
  assign n262 = n253 & n261 ;
  assign n263 = ( n236 & n259 ) | ( n236 & n262 ) | ( n259 & n262 ) ;
  assign n264 = n260 | n263 ;
  assign n265 = n238 & n262 ;
  assign n266 = ( n216 & n264 ) | ( n216 & n265 ) | ( n264 & n265 ) ;
  assign n267 = n264 | n266 ;
  assign n269 = n268 ^ n267 ^ 1'b0 ;
  assign n271 = ( x24 & x88 ) | ( x24 & n267 ) | ( x88 & n267 ) ;
  assign n270 = x89 ^ x25 ^ 1'b0 ;
  assign n272 = n271 ^ n270 ^ 1'b0 ;
  assign n278 = x90 ^ x26 ^ 1'b0 ;
  assign n273 = x24 & x88 ;
  assign n274 = ( x25 & x89 ) | ( x25 & n273 ) | ( x89 & n273 ) ;
  assign n275 = n268 & n270 ;
  assign n276 = ( n267 & n274 ) | ( n267 & n275 ) | ( n274 & n275 ) ;
  assign n277 = n274 | n276 ;
  assign n279 = n278 ^ n277 ^ 1'b0 ;
  assign n281 = ( x26 & x90 ) | ( x26 & n277 ) | ( x90 & n277 ) ;
  assign n280 = x91 ^ x27 ^ 1'b0 ;
  assign n282 = n281 ^ n280 ^ 1'b0 ;
  assign n292 = x92 ^ x28 ^ 1'b0 ;
  assign n283 = x26 & x90 ;
  assign n284 = ( x27 & x91 ) | ( x27 & n283 ) | ( x91 & n283 ) ;
  assign n285 = n278 & n280 ;
  assign n286 = ( n274 & n284 ) | ( n274 & n285 ) | ( n284 & n285 ) ;
  assign n287 = n284 | n286 ;
  assign n288 = ( n275 & n278 ) | ( n275 & ~n280 ) | ( n278 & ~n280 ) ;
  assign n289 = n280 & n288 ;
  assign n290 = ( n267 & n287 ) | ( n267 & n289 ) | ( n287 & n289 ) ;
  assign n291 = n287 | n290 ;
  assign n293 = n292 ^ n291 ^ 1'b0 ;
  assign n295 = ( x28 & x92 ) | ( x28 & n291 ) | ( x92 & n291 ) ;
  assign n294 = x93 ^ x29 ^ 1'b0 ;
  assign n296 = n295 ^ n294 ^ 1'b0 ;
  assign n302 = x94 ^ x30 ^ 1'b0 ;
  assign n297 = x28 & x92 ;
  assign n298 = ( x29 & x93 ) | ( x29 & n297 ) | ( x93 & n297 ) ;
  assign n299 = n292 & n294 ;
  assign n300 = ( n291 & n298 ) | ( n291 & n299 ) | ( n298 & n299 ) ;
  assign n301 = n298 | n300 ;
  assign n303 = n302 ^ n301 ^ 1'b0 ;
  assign n305 = ( x30 & x94 ) | ( x30 & n301 ) | ( x94 & n301 ) ;
  assign n304 = x95 ^ x31 ^ 1'b0 ;
  assign n306 = n305 ^ n304 ^ 1'b0 ;
  assign n322 = x96 ^ x32 ^ 1'b0 ;
  assign n307 = x30 & x94 ;
  assign n308 = ( x31 & x95 ) | ( x31 & n307 ) | ( x95 & n307 ) ;
  assign n309 = ( n298 & n302 ) | ( n298 & ~n304 ) | ( n302 & ~n304 ) ;
  assign n310 = n304 & n309 ;
  assign n311 = n308 | n310 ;
  assign n312 = ( n299 & n302 ) | ( n299 & ~n304 ) | ( n302 & ~n304 ) ;
  assign n313 = n304 & n312 ;
  assign n314 = ( n287 & n310 ) | ( n287 & n313 ) | ( n310 & n313 ) ;
  assign n315 = n311 | n314 ;
  assign n316 = n289 & n313 ;
  assign n317 = ( n264 & n315 ) | ( n264 & n316 ) | ( n315 & n316 ) ;
  assign n318 = n315 | n317 ;
  assign n319 = ~n216 & n265 ;
  assign n320 = ( n265 & n316 ) | ( n265 & n319 ) | ( n316 & n319 ) ;
  assign n321 = ( n318 & ~n319 ) | ( n318 & n320 ) | ( ~n319 & n320 ) ;
  assign n323 = n322 ^ n321 ^ 1'b0 ;
  assign n325 = ( x32 & x96 ) | ( x32 & n321 ) | ( x96 & n321 ) ;
  assign n324 = x97 ^ x33 ^ 1'b0 ;
  assign n326 = n325 ^ n324 ^ 1'b0 ;
  assign n332 = x98 ^ x34 ^ 1'b0 ;
  assign n327 = x32 & x96 ;
  assign n328 = ( x33 & x97 ) | ( x33 & n327 ) | ( x97 & n327 ) ;
  assign n329 = n322 & n324 ;
  assign n330 = ( n321 & n328 ) | ( n321 & n329 ) | ( n328 & n329 ) ;
  assign n331 = n328 | n330 ;
  assign n333 = n332 ^ n331 ^ 1'b0 ;
  assign n335 = ( x34 & x98 ) | ( x34 & n331 ) | ( x98 & n331 ) ;
  assign n334 = x99 ^ x35 ^ 1'b0 ;
  assign n336 = n335 ^ n334 ^ 1'b0 ;
  assign n346 = x100 ^ x36 ^ 1'b0 ;
  assign n337 = x34 & x98 ;
  assign n338 = ( x35 & x99 ) | ( x35 & n337 ) | ( x99 & n337 ) ;
  assign n339 = n332 & n334 ;
  assign n340 = ( n328 & n338 ) | ( n328 & n339 ) | ( n338 & n339 ) ;
  assign n341 = n338 | n340 ;
  assign n342 = ( n329 & n332 ) | ( n329 & ~n334 ) | ( n332 & ~n334 ) ;
  assign n343 = n334 & n342 ;
  assign n344 = ( n321 & n341 ) | ( n321 & n343 ) | ( n341 & n343 ) ;
  assign n345 = n341 | n344 ;
  assign n347 = n346 ^ n345 ^ 1'b0 ;
  assign n349 = ( x36 & x100 ) | ( x36 & n345 ) | ( x100 & n345 ) ;
  assign n348 = x101 ^ x37 ^ 1'b0 ;
  assign n350 = n349 ^ n348 ^ 1'b0 ;
  assign n356 = x102 ^ x38 ^ 1'b0 ;
  assign n351 = x36 & x100 ;
  assign n352 = ( x37 & x101 ) | ( x37 & n351 ) | ( x101 & n351 ) ;
  assign n353 = n346 & n348 ;
  assign n354 = ( n345 & n352 ) | ( n345 & n353 ) | ( n352 & n353 ) ;
  assign n355 = n352 | n354 ;
  assign n357 = n356 ^ n355 ^ 1'b0 ;
  assign n359 = ( x38 & x102 ) | ( x38 & n355 ) | ( x102 & n355 ) ;
  assign n358 = x103 ^ x39 ^ 1'b0 ;
  assign n360 = n359 ^ n358 ^ 1'b0 ;
  assign n373 = x104 ^ x40 ^ 1'b0 ;
  assign n361 = x38 & x102 ;
  assign n362 = ( x39 & x103 ) | ( x39 & n361 ) | ( x103 & n361 ) ;
  assign n363 = ( n352 & n356 ) | ( n352 & ~n358 ) | ( n356 & ~n358 ) ;
  assign n364 = n358 & n363 ;
  assign n365 = n362 | n364 ;
  assign n366 = ( n353 & n356 ) | ( n353 & ~n358 ) | ( n356 & ~n358 ) ;
  assign n367 = n358 & n366 ;
  assign n368 = ( n341 & n364 ) | ( n341 & n367 ) | ( n364 & n367 ) ;
  assign n369 = n365 | n368 ;
  assign n370 = n343 & n367 ;
  assign n371 = ( n321 & n369 ) | ( n321 & n370 ) | ( n369 & n370 ) ;
  assign n372 = n369 | n371 ;
  assign n374 = n373 ^ n372 ^ 1'b0 ;
  assign n376 = ( x40 & x104 ) | ( x40 & n372 ) | ( x104 & n372 ) ;
  assign n375 = x105 ^ x41 ^ 1'b0 ;
  assign n377 = n376 ^ n375 ^ 1'b0 ;
  assign n383 = x106 ^ x42 ^ 1'b0 ;
  assign n378 = x40 & x104 ;
  assign n379 = ( x41 & x105 ) | ( x41 & n378 ) | ( x105 & n378 ) ;
  assign n380 = n373 & n375 ;
  assign n381 = ( n372 & n379 ) | ( n372 & n380 ) | ( n379 & n380 ) ;
  assign n382 = n379 | n381 ;
  assign n384 = n383 ^ n382 ^ 1'b0 ;
  assign n386 = ( x42 & x106 ) | ( x42 & n382 ) | ( x106 & n382 ) ;
  assign n385 = x107 ^ x43 ^ 1'b0 ;
  assign n387 = n386 ^ n385 ^ 1'b0 ;
  assign n397 = x108 ^ x44 ^ 1'b0 ;
  assign n388 = x42 & x106 ;
  assign n389 = ( x43 & x107 ) | ( x43 & n388 ) | ( x107 & n388 ) ;
  assign n390 = n383 & n385 ;
  assign n391 = ( n379 & n389 ) | ( n379 & n390 ) | ( n389 & n390 ) ;
  assign n392 = n389 | n391 ;
  assign n393 = ( n380 & n383 ) | ( n380 & ~n385 ) | ( n383 & ~n385 ) ;
  assign n394 = n385 & n393 ;
  assign n395 = ( n372 & n392 ) | ( n372 & n394 ) | ( n392 & n394 ) ;
  assign n396 = n392 | n395 ;
  assign n398 = n397 ^ n396 ^ 1'b0 ;
  assign n400 = ( x44 & x108 ) | ( x44 & n396 ) | ( x108 & n396 ) ;
  assign n399 = x109 ^ x45 ^ 1'b0 ;
  assign n401 = n400 ^ n399 ^ 1'b0 ;
  assign n407 = x110 ^ x46 ^ 1'b0 ;
  assign n402 = x44 & x108 ;
  assign n403 = ( x45 & x109 ) | ( x45 & n402 ) | ( x109 & n402 ) ;
  assign n404 = n397 & n399 ;
  assign n405 = ( n396 & n403 ) | ( n396 & n404 ) | ( n403 & n404 ) ;
  assign n406 = n403 | n405 ;
  assign n408 = n407 ^ n406 ^ 1'b0 ;
  assign n410 = ( x46 & x110 ) | ( x46 & n406 ) | ( x110 & n406 ) ;
  assign n409 = x111 ^ x47 ^ 1'b0 ;
  assign n411 = n410 ^ n409 ^ 1'b0 ;
  assign n427 = x112 ^ x48 ^ 1'b0 ;
  assign n412 = x46 & x110 ;
  assign n413 = ( x47 & x111 ) | ( x47 & n412 ) | ( x111 & n412 ) ;
  assign n414 = ( n403 & n407 ) | ( n403 & ~n409 ) | ( n407 & ~n409 ) ;
  assign n415 = n409 & n414 ;
  assign n416 = n413 | n415 ;
  assign n417 = ( n404 & n407 ) | ( n404 & ~n409 ) | ( n407 & ~n409 ) ;
  assign n418 = n409 & n417 ;
  assign n419 = ( n392 & n415 ) | ( n392 & n418 ) | ( n415 & n418 ) ;
  assign n420 = n416 | n419 ;
  assign n421 = n394 & n418 ;
  assign n422 = ( n369 & n420 ) | ( n369 & n421 ) | ( n420 & n421 ) ;
  assign n423 = n420 | n422 ;
  assign n424 = ~n321 & n370 ;
  assign n425 = ( n370 & n421 ) | ( n370 & n424 ) | ( n421 & n424 ) ;
  assign n426 = ( n423 & ~n424 ) | ( n423 & n425 ) | ( ~n424 & n425 ) ;
  assign n428 = n427 ^ n426 ^ 1'b0 ;
  assign n430 = ( x48 & x112 ) | ( x48 & n426 ) | ( x112 & n426 ) ;
  assign n429 = x113 ^ x49 ^ 1'b0 ;
  assign n431 = n430 ^ n429 ^ 1'b0 ;
  assign n437 = x114 ^ x50 ^ 1'b0 ;
  assign n432 = x48 & x112 ;
  assign n433 = ( x49 & x113 ) | ( x49 & n432 ) | ( x113 & n432 ) ;
  assign n434 = n427 & n429 ;
  assign n435 = ( n426 & n433 ) | ( n426 & n434 ) | ( n433 & n434 ) ;
  assign n436 = n433 | n435 ;
  assign n438 = n437 ^ n436 ^ 1'b0 ;
  assign n440 = ( x50 & x114 ) | ( x50 & n436 ) | ( x114 & n436 ) ;
  assign n439 = x115 ^ x51 ^ 1'b0 ;
  assign n441 = n440 ^ n439 ^ 1'b0 ;
  assign n451 = x116 ^ x52 ^ 1'b0 ;
  assign n442 = x50 & x114 ;
  assign n443 = ( x51 & x115 ) | ( x51 & n442 ) | ( x115 & n442 ) ;
  assign n444 = n437 & n439 ;
  assign n445 = ( n433 & n443 ) | ( n433 & n444 ) | ( n443 & n444 ) ;
  assign n446 = n443 | n445 ;
  assign n447 = ( n434 & n437 ) | ( n434 & ~n439 ) | ( n437 & ~n439 ) ;
  assign n448 = n439 & n447 ;
  assign n449 = ( n426 & n446 ) | ( n426 & n448 ) | ( n446 & n448 ) ;
  assign n450 = n446 | n449 ;
  assign n452 = n451 ^ n450 ^ 1'b0 ;
  assign n454 = ( x52 & x116 ) | ( x52 & n450 ) | ( x116 & n450 ) ;
  assign n453 = x117 ^ x53 ^ 1'b0 ;
  assign n455 = n454 ^ n453 ^ 1'b0 ;
  assign n461 = x118 ^ x54 ^ 1'b0 ;
  assign n456 = x52 & x116 ;
  assign n457 = ( x53 & x117 ) | ( x53 & n456 ) | ( x117 & n456 ) ;
  assign n458 = n451 & n453 ;
  assign n459 = ( n450 & n457 ) | ( n450 & n458 ) | ( n457 & n458 ) ;
  assign n460 = n457 | n459 ;
  assign n462 = n461 ^ n460 ^ 1'b0 ;
  assign n464 = ( x54 & x118 ) | ( x54 & n460 ) | ( x118 & n460 ) ;
  assign n463 = x119 ^ x55 ^ 1'b0 ;
  assign n465 = n464 ^ n463 ^ 1'b0 ;
  assign n478 = x120 ^ x56 ^ 1'b0 ;
  assign n466 = x54 & x118 ;
  assign n467 = ( x55 & x119 ) | ( x55 & n466 ) | ( x119 & n466 ) ;
  assign n468 = ( n457 & n461 ) | ( n457 & ~n463 ) | ( n461 & ~n463 ) ;
  assign n469 = n463 & n468 ;
  assign n470 = n467 | n469 ;
  assign n471 = ( n458 & n461 ) | ( n458 & ~n463 ) | ( n461 & ~n463 ) ;
  assign n472 = n463 & n471 ;
  assign n473 = ( n446 & n469 ) | ( n446 & n472 ) | ( n469 & n472 ) ;
  assign n474 = n470 | n473 ;
  assign n475 = ~n426 & n448 ;
  assign n476 = ( n448 & n472 ) | ( n448 & n475 ) | ( n472 & n475 ) ;
  assign n477 = ( n474 & ~n475 ) | ( n474 & n476 ) | ( ~n475 & n476 ) ;
  assign n479 = n478 ^ n477 ^ 1'b0 ;
  assign n481 = ( x56 & x120 ) | ( x56 & n477 ) | ( x120 & n477 ) ;
  assign n480 = x121 ^ x57 ^ 1'b0 ;
  assign n482 = n481 ^ n480 ^ 1'b0 ;
  assign n488 = x122 ^ x58 ^ 1'b0 ;
  assign n483 = x56 & x120 ;
  assign n484 = ( x57 & x121 ) | ( x57 & n483 ) | ( x121 & n483 ) ;
  assign n485 = n478 & n480 ;
  assign n486 = ( n477 & n484 ) | ( n477 & n485 ) | ( n484 & n485 ) ;
  assign n487 = n484 | n486 ;
  assign n489 = n488 ^ n487 ^ 1'b0 ;
  assign n491 = ( x58 & x122 ) | ( x58 & n487 ) | ( x122 & n487 ) ;
  assign n490 = x123 ^ x59 ^ 1'b0 ;
  assign n492 = n491 ^ n490 ^ 1'b0 ;
  assign n501 = x124 ^ x60 ^ 1'b0 ;
  assign n493 = x58 & x122 ;
  assign n494 = ( x59 & x123 ) | ( x59 & n493 ) | ( x123 & n493 ) ;
  assign n495 = n488 & n490 ;
  assign n496 = ( n484 & n494 ) | ( n484 & n495 ) | ( n494 & n495 ) ;
  assign n497 = n494 | n496 ;
  assign n498 = ~n477 & n485 ;
  assign n499 = ( n485 & n495 ) | ( n485 & n498 ) | ( n495 & n498 ) ;
  assign n500 = ( n497 & ~n498 ) | ( n497 & n499 ) | ( ~n498 & n499 ) ;
  assign n502 = n501 ^ n500 ^ 1'b0 ;
  assign n504 = ( x60 & x124 ) | ( x60 & n500 ) | ( x124 & n500 ) ;
  assign n503 = x125 ^ x61 ^ 1'b0 ;
  assign n505 = n504 ^ n503 ^ 1'b0 ;
  assign n511 = x126 ^ x62 ^ 1'b0 ;
  assign n506 = x60 & x124 ;
  assign n507 = ( x61 & x125 ) | ( x61 & n506 ) | ( x125 & n506 ) ;
  assign n508 = n500 & ~n501 ;
  assign n509 = ( n500 & n503 ) | ( n500 & n508 ) | ( n503 & n508 ) ;
  assign n510 = ( n507 & ~n508 ) | ( n507 & n509 ) | ( ~n508 & n509 ) ;
  assign n512 = n511 ^ n510 ^ 1'b0 ;
  assign n514 = ( x62 & x126 ) | ( x62 & n510 ) | ( x126 & n510 ) ;
  assign n513 = x127 ^ x63 ^ 1'b0 ;
  assign n515 = n514 ^ n513 ^ 1'b0 ;
  assign y0 = n129 ;
  assign y1 = n131 ;
  assign y2 = n134 ;
  assign y3 = n137 ;
  assign y4 = n144 ;
  assign y5 = n147 ;
  assign y6 = n154 ;
  assign y7 = n157 ;
  assign y8 = n167 ;
  assign y9 = n170 ;
  assign y10 = n177 ;
  assign y11 = n180 ;
  assign y12 = n191 ;
  assign y13 = n194 ;
  assign y14 = n201 ;
  assign y15 = n204 ;
  assign y16 = n218 ;
  assign y17 = n221 ;
  assign y18 = n228 ;
  assign y19 = n231 ;
  assign y20 = n242 ;
  assign y21 = n245 ;
  assign y22 = n252 ;
  assign y23 = n255 ;
  assign y24 = n269 ;
  assign y25 = n272 ;
  assign y26 = n279 ;
  assign y27 = n282 ;
  assign y28 = n293 ;
  assign y29 = n296 ;
  assign y30 = n303 ;
  assign y31 = n306 ;
  assign y32 = n323 ;
  assign y33 = n326 ;
  assign y34 = n333 ;
  assign y35 = n336 ;
  assign y36 = n347 ;
  assign y37 = n350 ;
  assign y38 = n357 ;
  assign y39 = n360 ;
  assign y40 = n374 ;
  assign y41 = n377 ;
  assign y42 = n384 ;
  assign y43 = n387 ;
  assign y44 = n398 ;
  assign y45 = n401 ;
  assign y46 = n408 ;
  assign y47 = n411 ;
  assign y48 = n428 ;
  assign y49 = n431 ;
  assign y50 = n438 ;
  assign y51 = n441 ;
  assign y52 = n452 ;
  assign y53 = n455 ;
  assign y54 = n462 ;
  assign y55 = n465 ;
  assign y56 = n479 ;
  assign y57 = n482 ;
  assign y58 = n489 ;
  assign y59 = n492 ;
  assign y60 = n502 ;
  assign y61 = n505 ;
  assign y62 = n512 ;
  assign y63 = n515 ;
endmodule
