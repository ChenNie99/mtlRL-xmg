module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 ;
  assign n129 = x64 ^ x0 ^ 1'b0 ;
  assign n130 = x0 & x64 ;
  assign n131 = n130 ^ x65 ^ x1 ;
  assign n133 = ( x1 & x65 ) | ( x1 & n130 ) | ( x65 & n130 ) ;
  assign n132 = x66 ^ x2 ^ 1'b0 ;
  assign n134 = n133 ^ n132 ^ 1'b0 ;
  assign n136 = ( x2 & x66 ) | ( x2 & n133 ) | ( x66 & n133 ) ;
  assign n135 = x67 ^ x3 ^ 1'b0 ;
  assign n137 = n136 ^ n135 ^ 1'b0 ;
  assign n139 = x2 & x66 ;
  assign n140 = ( x3 & x67 ) | ( x3 & n139 ) | ( x67 & n139 ) ;
  assign n141 = n132 & n135 ;
  assign n142 = ( n133 & n140 ) | ( n133 & n141 ) | ( n140 & n141 ) ;
  assign n143 = n140 | n142 ;
  assign n138 = x68 ^ x4 ^ 1'b0 ;
  assign n144 = n143 ^ n138 ^ 1'b0 ;
  assign n146 = ( x4 & x68 ) | ( x4 & n143 ) | ( x68 & n143 ) ;
  assign n145 = x69 ^ x5 ^ 1'b0 ;
  assign n147 = n146 ^ n145 ^ 1'b0 ;
  assign n149 = x4 & x68 ;
  assign n150 = ( x5 & x69 ) | ( x5 & n149 ) | ( x69 & n149 ) ;
  assign n151 = n138 & n145 ;
  assign n152 = ( n143 & n150 ) | ( n143 & n151 ) | ( n150 & n151 ) ;
  assign n153 = n150 | n152 ;
  assign n148 = x70 ^ x6 ^ 1'b0 ;
  assign n154 = n153 ^ n148 ^ 1'b0 ;
  assign n156 = ( x6 & x70 ) | ( x6 & n153 ) | ( x70 & n153 ) ;
  assign n155 = x71 ^ x7 ^ 1'b0 ;
  assign n157 = n156 ^ n155 ^ 1'b0 ;
  assign n159 = x6 & x70 ;
  assign n160 = ( x7 & x71 ) | ( x7 & n159 ) | ( x71 & n159 ) ;
  assign n161 = n148 & n155 ;
  assign n162 = n143 & n151 ;
  assign n163 = n161 & n162 ;
  assign n164 = n150 & n161 ;
  assign n165 = n163 | n164 ;
  assign n166 = n160 | n165 ;
  assign n158 = x72 ^ x8 ^ 1'b0 ;
  assign n167 = n166 ^ n158 ^ 1'b0 ;
  assign n169 = ( x8 & x72 ) | ( x8 & n166 ) | ( x72 & n166 ) ;
  assign n168 = x73 ^ x9 ^ 1'b0 ;
  assign n170 = n169 ^ n168 ^ 1'b0 ;
  assign n172 = x8 & x72 ;
  assign n173 = ( x9 & x73 ) | ( x9 & n172 ) | ( x73 & n172 ) ;
  assign n174 = n158 & n168 ;
  assign n175 = ( n166 & n173 ) | ( n166 & n174 ) | ( n173 & n174 ) ;
  assign n176 = n173 | n175 ;
  assign n171 = x74 ^ x10 ^ 1'b0 ;
  assign n177 = n176 ^ n171 ^ 1'b0 ;
  assign n179 = ( x10 & x74 ) | ( x10 & n176 ) | ( x74 & n176 ) ;
  assign n178 = x75 ^ x11 ^ 1'b0 ;
  assign n180 = n179 ^ n178 ^ 1'b0 ;
  assign n182 = x10 & x74 ;
  assign n183 = ( x11 & x75 ) | ( x11 & n182 ) | ( x75 & n182 ) ;
  assign n184 = n171 & n178 ;
  assign n185 = ( n173 & n183 ) | ( n173 & n184 ) | ( n183 & n184 ) ;
  assign n186 = n183 | n185 ;
  assign n187 = n174 & n184 ;
  assign n188 = ( n166 & n186 ) | ( n166 & n187 ) | ( n186 & n187 ) ;
  assign n189 = n186 | n188 ;
  assign n181 = x76 ^ x12 ^ 1'b0 ;
  assign n190 = n189 ^ n181 ^ 1'b0 ;
  assign n192 = ( x12 & x76 ) | ( x12 & n189 ) | ( x76 & n189 ) ;
  assign n191 = x77 ^ x13 ^ 1'b0 ;
  assign n193 = n192 ^ n191 ^ 1'b0 ;
  assign n195 = x12 & x76 ;
  assign n196 = ( x13 & x77 ) | ( x13 & n195 ) | ( x77 & n195 ) ;
  assign n197 = n181 & n191 ;
  assign n198 = ( n189 & n196 ) | ( n189 & n197 ) | ( n196 & n197 ) ;
  assign n199 = n196 | n198 ;
  assign n194 = x78 ^ x14 ^ 1'b0 ;
  assign n200 = n199 ^ n194 ^ 1'b0 ;
  assign n202 = ( x14 & x78 ) | ( x14 & n199 ) | ( x78 & n199 ) ;
  assign n201 = x79 ^ x15 ^ 1'b0 ;
  assign n203 = n202 ^ n201 ^ 1'b0 ;
  assign n205 = x14 & x78 ;
  assign n206 = ( x15 & x79 ) | ( x15 & n205 ) | ( x79 & n205 ) ;
  assign n207 = n194 & n201 ;
  assign n208 = n197 & n207 ;
  assign n209 = n186 & n208 ;
  assign n210 = n196 & n207 ;
  assign n211 = n209 | n210 ;
  assign n212 = n206 | n211 ;
  assign n213 = n187 & n208 ;
  assign n214 = ( n166 & n212 ) | ( n166 & n213 ) | ( n212 & n213 ) ;
  assign n215 = n212 | n214 ;
  assign n204 = x80 ^ x16 ^ 1'b0 ;
  assign n216 = n215 ^ n204 ^ 1'b0 ;
  assign n218 = ( x16 & x80 ) | ( x16 & n215 ) | ( x80 & n215 ) ;
  assign n217 = x81 ^ x17 ^ 1'b0 ;
  assign n219 = n218 ^ n217 ^ 1'b0 ;
  assign n221 = x16 & x80 ;
  assign n222 = ( x17 & x81 ) | ( x17 & n221 ) | ( x81 & n221 ) ;
  assign n223 = n204 & n217 ;
  assign n224 = ( n215 & n222 ) | ( n215 & n223 ) | ( n222 & n223 ) ;
  assign n225 = n222 | n224 ;
  assign n220 = x82 ^ x18 ^ 1'b0 ;
  assign n226 = n225 ^ n220 ^ 1'b0 ;
  assign n228 = ( x18 & x82 ) | ( x18 & n225 ) | ( x82 & n225 ) ;
  assign n227 = x83 ^ x19 ^ 1'b0 ;
  assign n229 = n228 ^ n227 ^ 1'b0 ;
  assign n231 = x18 & x82 ;
  assign n232 = ( x19 & x83 ) | ( x19 & n231 ) | ( x83 & n231 ) ;
  assign n233 = n220 & n227 ;
  assign n234 = ( n222 & n232 ) | ( n222 & n233 ) | ( n232 & n233 ) ;
  assign n235 = n232 | n234 ;
  assign n236 = n223 & n233 ;
  assign n237 = ( n215 & n235 ) | ( n215 & n236 ) | ( n235 & n236 ) ;
  assign n238 = n235 | n237 ;
  assign n230 = x84 ^ x20 ^ 1'b0 ;
  assign n239 = n238 ^ n230 ^ 1'b0 ;
  assign n241 = ( x20 & x84 ) | ( x20 & n238 ) | ( x84 & n238 ) ;
  assign n240 = x85 ^ x21 ^ 1'b0 ;
  assign n242 = n241 ^ n240 ^ 1'b0 ;
  assign n244 = x20 & x84 ;
  assign n245 = ( x21 & x85 ) | ( x21 & n244 ) | ( x85 & n244 ) ;
  assign n246 = n230 & n240 ;
  assign n247 = ( n238 & n245 ) | ( n238 & n246 ) | ( n245 & n246 ) ;
  assign n248 = n245 | n247 ;
  assign n243 = x86 ^ x22 ^ 1'b0 ;
  assign n249 = n248 ^ n243 ^ 1'b0 ;
  assign n251 = ( x22 & x86 ) | ( x22 & n248 ) | ( x86 & n248 ) ;
  assign n250 = x87 ^ x23 ^ 1'b0 ;
  assign n252 = n251 ^ n250 ^ 1'b0 ;
  assign n254 = x22 & x86 ;
  assign n255 = ( x23 & x87 ) | ( x23 & n254 ) | ( x87 & n254 ) ;
  assign n256 = n243 & n250 ;
  assign n257 = n246 & n256 ;
  assign n258 = n235 & n257 ;
  assign n259 = n245 & n256 ;
  assign n260 = n258 | n259 ;
  assign n261 = n255 | n260 ;
  assign n262 = n236 & n257 ;
  assign n263 = ( n215 & n261 ) | ( n215 & n262 ) | ( n261 & n262 ) ;
  assign n264 = n261 | n263 ;
  assign n253 = x88 ^ x24 ^ 1'b0 ;
  assign n265 = n264 ^ n253 ^ 1'b0 ;
  assign n267 = ( x24 & x88 ) | ( x24 & n264 ) | ( x88 & n264 ) ;
  assign n266 = x89 ^ x25 ^ 1'b0 ;
  assign n268 = n267 ^ n266 ^ 1'b0 ;
  assign n270 = x24 & x88 ;
  assign n271 = ( x25 & x89 ) | ( x25 & n270 ) | ( x89 & n270 ) ;
  assign n272 = n253 & n266 ;
  assign n273 = ( n264 & n271 ) | ( n264 & n272 ) | ( n271 & n272 ) ;
  assign n274 = n271 | n273 ;
  assign n269 = x90 ^ x26 ^ 1'b0 ;
  assign n275 = n274 ^ n269 ^ 1'b0 ;
  assign n277 = ( x26 & x90 ) | ( x26 & n274 ) | ( x90 & n274 ) ;
  assign n276 = x91 ^ x27 ^ 1'b0 ;
  assign n278 = n277 ^ n276 ^ 1'b0 ;
  assign n280 = x26 & x90 ;
  assign n281 = ( x27 & x91 ) | ( x27 & n280 ) | ( x91 & n280 ) ;
  assign n282 = n269 & n276 ;
  assign n283 = ( n271 & n281 ) | ( n271 & n282 ) | ( n281 & n282 ) ;
  assign n284 = n281 | n283 ;
  assign n285 = n272 & n282 ;
  assign n286 = ( n264 & n284 ) | ( n264 & n285 ) | ( n284 & n285 ) ;
  assign n287 = n284 | n286 ;
  assign n279 = x92 ^ x28 ^ 1'b0 ;
  assign n288 = n287 ^ n279 ^ 1'b0 ;
  assign n290 = ( x28 & x92 ) | ( x28 & n287 ) | ( x92 & n287 ) ;
  assign n289 = x93 ^ x29 ^ 1'b0 ;
  assign n291 = n290 ^ n289 ^ 1'b0 ;
  assign n293 = x28 & x92 ;
  assign n294 = ( x29 & x93 ) | ( x29 & n293 ) | ( x93 & n293 ) ;
  assign n295 = n279 & n289 ;
  assign n296 = ( n287 & n294 ) | ( n287 & n295 ) | ( n294 & n295 ) ;
  assign n297 = n294 | n296 ;
  assign n292 = x94 ^ x30 ^ 1'b0 ;
  assign n298 = n297 ^ n292 ^ 1'b0 ;
  assign n300 = ( x30 & x94 ) | ( x30 & n297 ) | ( x94 & n297 ) ;
  assign n299 = x95 ^ x31 ^ 1'b0 ;
  assign n301 = n300 ^ n299 ^ 1'b0 ;
  assign n303 = x30 & x94 ;
  assign n304 = ( x31 & x95 ) | ( x31 & n303 ) | ( x95 & n303 ) ;
  assign n305 = n292 & n299 ;
  assign n306 = n295 & n305 ;
  assign n307 = n284 & n306 ;
  assign n308 = n294 & n305 ;
  assign n309 = n307 | n308 ;
  assign n310 = n304 | n309 ;
  assign n311 = n285 & n306 ;
  assign n312 = ( n261 & n310 ) | ( n261 & n311 ) | ( n310 & n311 ) ;
  assign n313 = n310 | n312 ;
  assign n314 = n262 & n311 ;
  assign n315 = ( n215 & n313 ) | ( n215 & n314 ) | ( n313 & n314 ) ;
  assign n316 = n313 | n315 ;
  assign n302 = x96 ^ x32 ^ 1'b0 ;
  assign n317 = n316 ^ n302 ^ 1'b0 ;
  assign n319 = ( x32 & x96 ) | ( x32 & n316 ) | ( x96 & n316 ) ;
  assign n318 = x97 ^ x33 ^ 1'b0 ;
  assign n320 = n319 ^ n318 ^ 1'b0 ;
  assign n322 = x32 & x96 ;
  assign n323 = ( x33 & x97 ) | ( x33 & n322 ) | ( x97 & n322 ) ;
  assign n324 = n302 & n318 ;
  assign n325 = ( n316 & n323 ) | ( n316 & n324 ) | ( n323 & n324 ) ;
  assign n326 = n323 | n325 ;
  assign n321 = x98 ^ x34 ^ 1'b0 ;
  assign n327 = n326 ^ n321 ^ 1'b0 ;
  assign n329 = ( x34 & x98 ) | ( x34 & n326 ) | ( x98 & n326 ) ;
  assign n328 = x99 ^ x35 ^ 1'b0 ;
  assign n330 = n329 ^ n328 ^ 1'b0 ;
  assign n332 = x34 & x98 ;
  assign n333 = ( x35 & x99 ) | ( x35 & n332 ) | ( x99 & n332 ) ;
  assign n334 = n321 & n328 ;
  assign n335 = ( n323 & n333 ) | ( n323 & n334 ) | ( n333 & n334 ) ;
  assign n336 = n333 | n335 ;
  assign n337 = n324 & n334 ;
  assign n338 = ( n316 & n336 ) | ( n316 & n337 ) | ( n336 & n337 ) ;
  assign n339 = n336 | n338 ;
  assign n331 = x100 ^ x36 ^ 1'b0 ;
  assign n340 = n339 ^ n331 ^ 1'b0 ;
  assign n342 = ( x36 & x100 ) | ( x36 & n339 ) | ( x100 & n339 ) ;
  assign n341 = x101 ^ x37 ^ 1'b0 ;
  assign n343 = n342 ^ n341 ^ 1'b0 ;
  assign n345 = x36 & x100 ;
  assign n346 = ( x37 & x101 ) | ( x37 & n345 ) | ( x101 & n345 ) ;
  assign n347 = n331 & n341 ;
  assign n348 = ( n339 & n346 ) | ( n339 & n347 ) | ( n346 & n347 ) ;
  assign n349 = n346 | n348 ;
  assign n344 = x102 ^ x38 ^ 1'b0 ;
  assign n350 = n349 ^ n344 ^ 1'b0 ;
  assign n352 = ( x38 & x102 ) | ( x38 & n349 ) | ( x102 & n349 ) ;
  assign n351 = x103 ^ x39 ^ 1'b0 ;
  assign n353 = n352 ^ n351 ^ 1'b0 ;
  assign n355 = x38 & x102 ;
  assign n356 = ( x39 & x103 ) | ( x39 & n355 ) | ( x103 & n355 ) ;
  assign n357 = n344 & n351 ;
  assign n358 = n347 & n357 ;
  assign n359 = n336 & n358 ;
  assign n360 = n346 & n357 ;
  assign n361 = n359 | n360 ;
  assign n362 = n356 | n361 ;
  assign n363 = n337 & n358 ;
  assign n364 = ( n316 & n362 ) | ( n316 & n363 ) | ( n362 & n363 ) ;
  assign n365 = n362 | n364 ;
  assign n354 = x104 ^ x40 ^ 1'b0 ;
  assign n366 = n365 ^ n354 ^ 1'b0 ;
  assign n368 = ( x40 & x104 ) | ( x40 & n365 ) | ( x104 & n365 ) ;
  assign n367 = x105 ^ x41 ^ 1'b0 ;
  assign n369 = n368 ^ n367 ^ 1'b0 ;
  assign n371 = x40 & x104 ;
  assign n372 = ( x41 & x105 ) | ( x41 & n371 ) | ( x105 & n371 ) ;
  assign n373 = n354 & n367 ;
  assign n374 = ( n365 & n372 ) | ( n365 & n373 ) | ( n372 & n373 ) ;
  assign n375 = n372 | n374 ;
  assign n370 = x106 ^ x42 ^ 1'b0 ;
  assign n376 = n375 ^ n370 ^ 1'b0 ;
  assign n378 = ( x42 & x106 ) | ( x42 & n375 ) | ( x106 & n375 ) ;
  assign n377 = x107 ^ x43 ^ 1'b0 ;
  assign n379 = n378 ^ n377 ^ 1'b0 ;
  assign n381 = x42 & x106 ;
  assign n382 = ( x43 & x107 ) | ( x43 & n381 ) | ( x107 & n381 ) ;
  assign n383 = n370 & n377 ;
  assign n384 = ( n372 & n382 ) | ( n372 & n383 ) | ( n382 & n383 ) ;
  assign n385 = n382 | n384 ;
  assign n386 = n373 & n383 ;
  assign n387 = ( n365 & n385 ) | ( n365 & n386 ) | ( n385 & n386 ) ;
  assign n388 = n385 | n387 ;
  assign n380 = x108 ^ x44 ^ 1'b0 ;
  assign n389 = n388 ^ n380 ^ 1'b0 ;
  assign n391 = ( x44 & x108 ) | ( x44 & n388 ) | ( x108 & n388 ) ;
  assign n390 = x109 ^ x45 ^ 1'b0 ;
  assign n392 = n391 ^ n390 ^ 1'b0 ;
  assign n394 = x44 & x108 ;
  assign n395 = ( x45 & x109 ) | ( x45 & n394 ) | ( x109 & n394 ) ;
  assign n396 = n380 & n390 ;
  assign n397 = ( n388 & n395 ) | ( n388 & n396 ) | ( n395 & n396 ) ;
  assign n398 = n395 | n397 ;
  assign n393 = x110 ^ x46 ^ 1'b0 ;
  assign n399 = n398 ^ n393 ^ 1'b0 ;
  assign n401 = ( x46 & x110 ) | ( x46 & n398 ) | ( x110 & n398 ) ;
  assign n400 = x111 ^ x47 ^ 1'b0 ;
  assign n402 = n401 ^ n400 ^ 1'b0 ;
  assign n404 = x46 & x110 ;
  assign n405 = ( x47 & x111 ) | ( x47 & n404 ) | ( x111 & n404 ) ;
  assign n406 = n393 & n400 ;
  assign n407 = n396 & n406 ;
  assign n408 = n385 & n407 ;
  assign n409 = n395 & n406 ;
  assign n410 = n408 | n409 ;
  assign n411 = n405 | n410 ;
  assign n412 = n386 & n407 ;
  assign n413 = ( n362 & n411 ) | ( n362 & n412 ) | ( n411 & n412 ) ;
  assign n414 = n411 | n413 ;
  assign n415 = n363 & n412 ;
  assign n416 = ( n316 & n414 ) | ( n316 & n415 ) | ( n414 & n415 ) ;
  assign n417 = n414 | n416 ;
  assign n403 = x112 ^ x48 ^ 1'b0 ;
  assign n418 = n417 ^ n403 ^ 1'b0 ;
  assign n420 = ( x48 & x112 ) | ( x48 & n417 ) | ( x112 & n417 ) ;
  assign n419 = x113 ^ x49 ^ 1'b0 ;
  assign n421 = n420 ^ n419 ^ 1'b0 ;
  assign n423 = x48 & x112 ;
  assign n424 = ( x49 & x113 ) | ( x49 & n423 ) | ( x113 & n423 ) ;
  assign n425 = n403 & n419 ;
  assign n426 = ( n417 & n424 ) | ( n417 & n425 ) | ( n424 & n425 ) ;
  assign n427 = n424 | n426 ;
  assign n422 = x114 ^ x50 ^ 1'b0 ;
  assign n428 = n427 ^ n422 ^ 1'b0 ;
  assign n430 = ( x50 & x114 ) | ( x50 & n427 ) | ( x114 & n427 ) ;
  assign n429 = x115 ^ x51 ^ 1'b0 ;
  assign n431 = n430 ^ n429 ^ 1'b0 ;
  assign n433 = x50 & x114 ;
  assign n434 = ( x51 & x115 ) | ( x51 & n433 ) | ( x115 & n433 ) ;
  assign n435 = n422 & n429 ;
  assign n436 = ( n424 & n434 ) | ( n424 & n435 ) | ( n434 & n435 ) ;
  assign n437 = n434 | n436 ;
  assign n438 = n425 & n435 ;
  assign n439 = ( n417 & n437 ) | ( n417 & n438 ) | ( n437 & n438 ) ;
  assign n440 = n437 | n439 ;
  assign n432 = x116 ^ x52 ^ 1'b0 ;
  assign n441 = n440 ^ n432 ^ 1'b0 ;
  assign n443 = ( x52 & x116 ) | ( x52 & n440 ) | ( x116 & n440 ) ;
  assign n442 = x117 ^ x53 ^ 1'b0 ;
  assign n444 = n443 ^ n442 ^ 1'b0 ;
  assign n446 = x52 & x116 ;
  assign n447 = ( x53 & x117 ) | ( x53 & n446 ) | ( x117 & n446 ) ;
  assign n448 = n432 & n442 ;
  assign n449 = ( n440 & n447 ) | ( n440 & n448 ) | ( n447 & n448 ) ;
  assign n450 = n447 | n449 ;
  assign n445 = x118 ^ x54 ^ 1'b0 ;
  assign n451 = n450 ^ n445 ^ 1'b0 ;
  assign n453 = ( x54 & x118 ) | ( x54 & n450 ) | ( x118 & n450 ) ;
  assign n452 = x119 ^ x55 ^ 1'b0 ;
  assign n454 = n453 ^ n452 ^ 1'b0 ;
  assign n456 = x54 & x118 ;
  assign n457 = ( x55 & x119 ) | ( x55 & n456 ) | ( x119 & n456 ) ;
  assign n458 = n445 & n452 ;
  assign n459 = n448 & n458 ;
  assign n460 = n437 & n459 ;
  assign n461 = n447 & n458 ;
  assign n462 = n460 | n461 ;
  assign n463 = n457 | n462 ;
  assign n464 = n438 & n459 ;
  assign n465 = ( n417 & n463 ) | ( n417 & n464 ) | ( n463 & n464 ) ;
  assign n466 = n463 | n465 ;
  assign n455 = x120 ^ x56 ^ 1'b0 ;
  assign n467 = n466 ^ n455 ^ 1'b0 ;
  assign n469 = ( x56 & x120 ) | ( x56 & n466 ) | ( x120 & n466 ) ;
  assign n468 = x121 ^ x57 ^ 1'b0 ;
  assign n470 = n469 ^ n468 ^ 1'b0 ;
  assign n472 = x56 & x120 ;
  assign n473 = ( x57 & x121 ) | ( x57 & n472 ) | ( x121 & n472 ) ;
  assign n474 = n455 & n468 ;
  assign n475 = ( n466 & n473 ) | ( n466 & n474 ) | ( n473 & n474 ) ;
  assign n476 = n473 | n475 ;
  assign n471 = x122 ^ x58 ^ 1'b0 ;
  assign n477 = n476 ^ n471 ^ 1'b0 ;
  assign n479 = ( x58 & x122 ) | ( x58 & n476 ) | ( x122 & n476 ) ;
  assign n478 = x123 ^ x59 ^ 1'b0 ;
  assign n480 = n479 ^ n478 ^ 1'b0 ;
  assign n482 = x58 & x122 ;
  assign n483 = ( x59 & x123 ) | ( x59 & n482 ) | ( x123 & n482 ) ;
  assign n484 = n471 & n478 ;
  assign n485 = n466 & n474 ;
  assign n486 = n484 & n485 ;
  assign n487 = n473 & n484 ;
  assign n488 = n486 | n487 ;
  assign n489 = n483 | n488 ;
  assign n481 = x124 ^ x60 ^ 1'b0 ;
  assign n490 = n489 ^ n481 ^ 1'b0 ;
  assign n492 = ( x60 & x124 ) | ( x60 & n489 ) | ( x124 & n489 ) ;
  assign n491 = x125 ^ x61 ^ 1'b0 ;
  assign n493 = n492 ^ n491 ^ 1'b0 ;
  assign n495 = x60 & x124 ;
  assign n496 = ( x61 & x125 ) | ( x61 & n495 ) | ( x125 & n495 ) ;
  assign n497 = n481 & n491 ;
  assign n498 = ( n489 & n496 ) | ( n489 & n497 ) | ( n496 & n497 ) ;
  assign n499 = n496 | n498 ;
  assign n494 = x126 ^ x62 ^ 1'b0 ;
  assign n500 = n499 ^ n494 ^ 1'b0 ;
  assign n502 = ( x62 & x126 ) | ( x62 & n499 ) | ( x126 & n499 ) ;
  assign n501 = x127 ^ x63 ^ 1'b0 ;
  assign n503 = n502 ^ n501 ^ 1'b0 ;
  assign y0 = n129 ;
  assign y1 = n131 ;
  assign y2 = n134 ;
  assign y3 = n137 ;
  assign y4 = n144 ;
  assign y5 = n147 ;
  assign y6 = n154 ;
  assign y7 = n157 ;
  assign y8 = n167 ;
  assign y9 = n170 ;
  assign y10 = n177 ;
  assign y11 = n180 ;
  assign y12 = n190 ;
  assign y13 = n193 ;
  assign y14 = n200 ;
  assign y15 = n203 ;
  assign y16 = n216 ;
  assign y17 = n219 ;
  assign y18 = n226 ;
  assign y19 = n229 ;
  assign y20 = n239 ;
  assign y21 = n242 ;
  assign y22 = n249 ;
  assign y23 = n252 ;
  assign y24 = n265 ;
  assign y25 = n268 ;
  assign y26 = n275 ;
  assign y27 = n278 ;
  assign y28 = n288 ;
  assign y29 = n291 ;
  assign y30 = n298 ;
  assign y31 = n301 ;
  assign y32 = n317 ;
  assign y33 = n320 ;
  assign y34 = n327 ;
  assign y35 = n330 ;
  assign y36 = n340 ;
  assign y37 = n343 ;
  assign y38 = n350 ;
  assign y39 = n353 ;
  assign y40 = n366 ;
  assign y41 = n369 ;
  assign y42 = n376 ;
  assign y43 = n379 ;
  assign y44 = n389 ;
  assign y45 = n392 ;
  assign y46 = n399 ;
  assign y47 = n402 ;
  assign y48 = n418 ;
  assign y49 = n421 ;
  assign y50 = n428 ;
  assign y51 = n431 ;
  assign y52 = n441 ;
  assign y53 = n444 ;
  assign y54 = n451 ;
  assign y55 = n454 ;
  assign y56 = n467 ;
  assign y57 = n470 ;
  assign y58 = n477 ;
  assign y59 = n480 ;
  assign y60 = n490 ;
  assign y61 = n493 ;
  assign y62 = n500 ;
  assign y63 = n503 ;
endmodule
